---------------------------------------------------------------------------------------------
--! @file   direct_mapped_ICache_tb.vhd
--! @author Nicolas Ruiz Requejo
--!
--! @Copyright  SPDX-FileCopyrightText: 2020 Nicolas Ruiz Requejo nicolas.r.requejo@gmail.com
--!             SPDX-License-Identifier: CERN-OHL-S-2.0+
--!
--!             This source is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,
--!             INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A
--!             PARTICULAR PURPOSE. Please see the CERN-OHL-S v2 for applicable conditions.
--!
--!             Source location: https://github.com/nicruireq/PeRISCore32
--!
--!             As per CERN-OHL-S v2 section 4, should You produce hardware based on this
--!             source, You must where practicable maintain the Source Location visible
--!             on the external case and documentation of the PeRISCore32 or other products 
--!             you make using this source.
--!
---------------------------------------------------------------------------------------------

-- VHDL Testbench Template 
-- Autogenerated from nicruireq::hdltools app 
-- Written by Nicolas Ruiz Requejo
-- 
-- Notice:
-- Fill this template with your test code
-- Please if you discover a bug submit an Issue in
-- https://github.com/nicruireq/XilinxTclStore
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.all;

library periscore32;
use periscore32.cpu_types.all;
use periscore32.testbench_helpers.all;

ENTITY direct_mapped_ICache_tb IS
END direct_mapped_ICache_tb;

ARCHITECTURE behavior OF direct_mapped_ICache_tb IS 

	-- Component Declaration for the Unit Under Test (UUT)
component direct_mapped_ICache is
    generic(
        address_bits : integer := 32; --! width in bits of input address
        index_width : integer := 8; --! number of lines of cache index
        block_size : integer := 32; --! size of cache block
        byte_select : integer := 2 --! number of bits to select byte in each block
    );
    port (
        clk : in std_logic;
        --enable : in std_logic;
        write_enable : in std_logic;
        --read_enable : in std_logic;
        address : in word;
        data_in : in word;
        data_out : out word
        --hit_miss : out std_logic
    );
end component;

	-- Inputs and Outputs
	signal clk : std_logic;
	signal write_enable : std_logic;
	signal address : word;
	signal data_in : word;
	signal data_out : word;

    constant clock_period: time := 10 ns;
    signal stop_the_clock: boolean;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	-- UUT:
	my_direct_mapped_icache : direct_mapped_ICache
	port map(
		clk => clk ,
		--enable => --enable ,
		write_enable => write_enable ,
		--read_enable => --read_enable ,
		address => address ,
		data_in => data_in ,
		data_out => data_out );

    clocking: process
    begin
        while not stop_the_clock loop
            clk <= '0', '1' after clock_period / 2;
            wait for clock_period;
        end loop;
        wait;
    end process;

   -- Stimulus process
   stim_proc: process
        variable addr_mod4 : 
            unsigned(address'length-1 downto 0) := x"00000000";
   begin

        -- Put initialisation code here
        wait for 20 ns;
	    -- Put test bench stimulus code here
        -- Writing
        write_enable <= '1';
        data_in <= rand_slv(data_in'length);
        address <= std_logic_vector(addr_mod4);
        wait for 10 ns;
        gen_address : while addr_mod4 < x"000003fc" loop
            addr_mod4 := addr_mod4 + x"00000004";
            address <= std_logic_vector(addr_mod4);
            data_in <= rand_slv(data_in'length);
            wait for 10 ns;
        end loop ; -- gen_address
        
        -- reading
        write_enable <= '0';
        address <= x"00000000";
        addr_mod4 := x"00000000";
        wait for 10 ns;
        while addr_mod4 < x"000003fc" loop
            addr_mod4 := addr_mod4 + x"00000004";
            address <= std_logic_vector(addr_mod4);
            wait for 10 ns;
        end loop ; 

        wait;
   end process;

END;
