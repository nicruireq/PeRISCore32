---------------------------------------------------------------------------------------------
--! @file   cpu_components.vhd
--! @author Nicolas Ruiz Requejo
--!
--! @Copyright  SPDX-FileCopyrightText: 2020 Nicolas Ruiz Requejo nicolas.r.requejo@gmail.com
--!             SPDX-License-Identifier: CERN-OHL-S-2.0+
--!
--!             This source is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,
--!             INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A
--!             PARTICULAR PURPOSE. Please see the CERN-OHL-S v2 for applicable conditions.
--!
--!             Source location: https://github.com/nicruireq/PeRISCore32
--!
--!             As per CERN-OHL-S v2 section 4, should You produce hardware based on this
--!             source, You must where practicable maintain the Source Location visible
--!             on the external case and documentation of the PeRISCore32 or other products 
--!             you make using this source.
--!
---------------------------------------------------------------------------------------------

-- VHDL Testbench Template 
-- Autogenerated from nicruireq::hdltools app 
-- Written by Nicolas Ruiz Requejo
-- 
-- Notice:
-- Fill this template with your test code
-- Please if you discover a bug submit an Issue in
-- https://github.com/nicruireq/XilinxTclStore
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

library periscore32;
use periscore32.cpu_types.all;
use periscore32.testbench_helpers.all;

ENTITY alu_tb IS
END alu_tb;

ARCHITECTURE behavior OF alu_tb IS 

	-- Component Declaration for the Unit Under Test (UUT)
component alu is
    generic (
        data_width : integer := 32;
        alu_control_width : integer := 5
    );
    port (
        operand_A : in std_logic_vector(data_width-1 downto 0);
        operand_B : in std_logic_vector(data_width-1 downto 0);
        control : in std_logic_vector(alu_control_width-1 downto 0);
        computation_out : out std_logic_vector(data_width-1 downto 0);
        zero_flag : out std_logic;
        overflow_flag : out std_logic
    ) ;
end component;
    
    constant data_width : integer := 32;
    constant alu_control_width : integer := 5;
	-- Inputs and Outputs
	signal operand_A : std_logic_vector(data_width-1 downto 0);
	signal operand_B : std_logic_vector(data_width-1 downto 0);
	signal control : std_logic_vector(alu_control_width-1 downto 0);
	signal computation_out : std_logic_vector(data_width-1 downto 0);
	signal zero_flag : std_logic;
	signal overflow_flag : std_logic;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	-- UUT:
	my_alu : alu
	generic map(
		data_width => 32,
		alu_control_width => 5)
	port map(
		operand_A => operand_A ,
		operand_B => operand_B ,
		control => control ,
		computation_out => computation_out ,
		zero_flag => zero_flag ,
		overflow_flag => overflow_flag );

   -- Stimulus process
   stim_proc: process
   begin
		-- two positive operands
		operand_A <= x"00001388";	-- 5000
		operand_B <= x"0008ff56";	-- 589654

		control <= alu_add;
		--wait for 50 ns;
		--assert computation_out = x"000912de" report "alu_add: bad result";
		--wait for 50 ns;
		assert_comb_eq(
			computation_out, x"000912de",
			"alu_add: bad result", 100 ns
		);

		control <= alu_add_unsigned;
		assert_comb_eq(
			computation_out, x"000912de",
			"alu_add_unsigned: bad result", 100 ns
		);
		--assert computation_out = x"000912de" report "alu_add_unsigned: bad result";
		--wait for 100 ns;

		control <= alu_sub;
		assert_comb_eq(
			computation_out, x"fff71432",
			"alu_sub: bad result", 100 ns
		);
		--assert computation_out = x"fff71432" report "alu_sub: bad result";
		--wait for 100 ns;

		control <= alu_sub_unsigned;
		assert_comb_eq(
			computation_out, x"fff71432",
			"alu_sub_unsigned: bad result",
			100 ns
		);
		--assert computation_out = x"fff71432" report "alu_sub_unsigned: bad result";
		--wait for 100 ns;

		control <= alu_set_on_less;
		assert_comb_eq(
			computation_out, x"00000001",
			"alu_set_on_less: bad result",
			100 ns
		);
		--assert computation_out = x"00000001" report "alu_set_on_less: bad result";
		--wait for 100 ns;

		control <= alu_set_on_less_unsigned;
		assert_comb_eq(
			computation_out, x"00000001",
			"alu_set_on_less_unsigned: bad result",
			100 ns
		);
		--assert computation_out = x"00000001" report "alu_set_on_less_unsigned: bad result";
		--wait for 100 ns;

		control <= alu_and;
		assert_comb_eq(
			computation_out, x"00001300",
			"alu_and: bad result", 100 ns
		);
		--assert computation_out = x"00001300" report "alu_and: bad result";
		--wait for 100 ns;

		control <= alu_xor;
		assert_comb_eq(
			computation_out, x"0008ecde",
			"alu_xor: bad result", 100 ns
		);
		--assert computation_out = x"0008ecde" report "alu_xor: bad result";
		--wait for 100 ns;

		control <= alu_nor;
		assert_comb_eq(
			computation_out, x"fff70021",
			"alu_nor: bad result", 100 ns
		);
		--assert computation_out = x"fff70021" report "alu_nor: bad result";
		--wait for 100 ns;
		
		control <= alu_or;
		assert_comb_eq(
			computation_out, x"0008ffde",
			"alu_or: bad result", 100 ns
		);
		--assert computation_out = x"0008ffde" report "alu_or: bad result";
		--wait for 100 ns;

		-- shifts with positive operand
		operand_A <= x"00000008";	-- 8
		operand_B <= x"00001388";	-- 5000
		control <= alu_sll;
		assert_comb_eq(
			computation_out, x"00138800",
			"alu_sll: bad result", 100 ns
		);
		--assert computation_out = x"00138800" report "alu_sll: bad result";
		--wait for 100 ns;

		control <= alu_slr;
		assert_comb_eq(
			computation_out, x"00000013",
			"alu_slr: bad result", 100 ns
		);
		--assert computation_out = x"00000013" report "alu_slr: bad result";
		--wait for 100 ns;

		control <= alu_sra;
		assert_comb_eq(
			computation_out, x"00000013",
			"alu_sra: bad result", 100 ns
		);
		--assert computation_out = x"00000013" report "alu_sra: bad result";
		--wait for 100 ns;

		-- shift right arithmetic with negative operand
		operand_B <= x"ff695b4c";	-- -9872564
		control <= alu_sra;
		assert_comb_eq(
			computation_out, x"ffff695b",
			"alu_sra: bad result", 100 ns
		);
		--assert computation_out = x"ffff695b" report "alu_sra: bad result";
		--wait for 100 ns;

		-- one negative and one positive
		operand_A <= x"ff695b4c";	-- -9872564
		operand_B <= x"0008ff56";
		control <= alu_add;
		assert_comb_eq(
			computation_out, x"ff725aa2",
			"alu_add: bad result", 100 ns
		);
		--assert computation_out = x"ff725aa2" report "alu_add: bad result";
		--wait for 100 ns;

		control <= alu_add_unsigned;
		assert_comb_eq(
			computation_out, x"ff725aa2",
			"alu_add_unsigned: bad result", 100 ns
		);
		--assert computation_out = x"ff725aa2" report "alu_add_unsigned: bad result";
		--wait for 100 ns;

		control <= alu_sub;
		assert_comb_eq(
			computation_out, x"ff605bf6",
			"alu_sub: bad result", 100 ns
		);
		--assert computation_out = x"ff605bf6" report "alu_sub: bad result";
		--wait for 100 ns;

		control <= alu_sub_unsigned;
		assert_comb_eq(
			computation_out, x"ff605bf6",
			"alu_sub_unsigned: bad result", 
			100 ns
		);
		--assert computation_out = x"ff605bf6" report "alu_sub_unsigned: bad result";
		--wait for 100 ns;

		control <= alu_set_on_less;
		assert_comb_eq(
			computation_out, x"00000001",
			"alu_set_on_less: bad result", 
			100 ns
		);
		--assert computation_out = x"00000001" report "alu_set_on_less: bad result";
		--wait for 100 ns;

		control <= alu_set_on_less_unsigned;
		assert_comb_eq(
			computation_out, x"00000000",
			"alu_set_on_less_unsigned: bad result", 
			100 ns
		);
		--assert computation_out = x"00000000" report "alu_set_on_less_unsigned: bad result";
		--wait for 100 ns;

		-- overflows testing
		operand_A <= x"80000000";
		operand_B <= x"ffffffff";
		
		control <= alu_add;
		assert_comb_eq(
			computation_out, x"7fffffff",
			"alu_add - signed add overflow result: bad", 
			100 ns
		);
		assert_comb_eq(
			overflow_flag, '1',
			"alu_add - signed add overflow not active", 
			0 ns
		);
		--assert computation_out = x"7fffffff" report "alu_add - signed add overflow result: bad";
		--assert overflow_flag = '1' report "alu_add - signed add overflow not active";
		--wait for 100 ns;

		control <= alu_add_unsigned;
		assert_comb_eq(
			computation_out, x"7fffffff",
			"alu_add_unsigned - unsigned add result: bad", 
			100 ns
		);
		assert_comb_eq(
			overflow_flag, '0',
			"alu_add_unsigned - unsigned add overflow must not be active", 
			0 ns
		);
		--assert computation_out = x"7fffffff" report "alu_add_unsigned - unsigned add result: bad";
		--assert overflow_flag = '0' report "alu_add_unsigned - unsigned add overflow must not be active";
		--wait for 100 ns;

		operand_B <= x"00000001";
		control <= alu_sub;
		assert_comb_eq(
			computation_out, x"7fffffff",
			"alu_sub - signed substract result: bad", 
			100 ns
		);
		assert_comb_eq(
			overflow_flag, '1',
			"alu_sub - signed substract overflow not active", 
			0 ns
		);
		--assert computation_out = x"7fffffff" report "alu_sub - signed substract result: bad";
		--assert overflow_flag = '1' report "alu_sub - signed substract overflow not active";
		--wait for 100 ns;

		control <= alu_sub_unsigned;
		assert_comb_eq(
			computation_out, x"7fffffff",
			"alu_sub_unsigned - unsigned substract result: bad", 
			100 ns
		);
		assert_comb_eq(
			overflow_flag, '0',
			"alu_sub_unsigned - unsigned substract overflow must not be active", 
			0 ns
		);
		--assert computation_out = x"7fffffff" report "alu_sub_unsigned - unsigned substract result: bad";
		--assert overflow_flag = '0' report "alu_sub_unsigned - unsigned substract overflow must not be active";
		--wait for 100 ns;

		-- lui, byte, half extensions
		operand_B <= x"00000819";
		control <= alu_lui;
		assert_comb_eq(
			computation_out, x"08190000",
			"alu_lui: bad result", 
			100 ns
		);
		--assert computation_out = x"08190000" report "alu_lui: bad result";
		--wait for 100 ns;

		control <= alu_extend_byte;
		assert_comb_eq(
			computation_out, x"00000019",
			"alu_extend_byte: positive byte bad result", 
			100 ns
		);
		--assert computation_out = x"00000019" report "alu_extend_byte: positive byte bad result";
		--wait for 100 ns;

		operand_B <= x"110010f7";
		control <= alu_extend_byte;
		assert_comb_eq(
			computation_out, x"fffffff7",
			"alu_extend_byte: negative byte bad result", 
			100 ns
		);
		--assert computation_out = x"fffffff7" report "alu_extend_byte: negative byte bad result";
		--wait for 100 ns;

		control <= alu_extend_half;
		assert_comb_eq(
			computation_out, x"000010f7",
			"alu_extend_half: positive halfword bad result", 
			100 ns
		);
		--assert computation_out = x"000010f7" report "alu_extend_half: positive halfword bad result";
		--wait for 100 ns;		
		
		operand_B <= x"0142ea60";	-- b15 to b0 -> -5536 
		control <= alu_extend_half;
		assert_comb_eq(
			computation_out, x"ffffea60",
			"alu_extend_half: negative halfword bad result", 
			100 ns
		);
		--assert computation_out = x"ffffea60" report "alu_extend_half: negative halfword bad result";
		--wait for 100 ns;

      wait;
   end process;

END;

